PACKAGE CommonLib IS

  function requiredBitNb (val : integer) return integer;

END CommonLib;
